module add_sub16(
    input [15:0] x,
    input [15:0] y,
    input cin,
    input sel,
    output [15:0] result,
    output cout, 
    output overflow
);
    

    wire
endmodule