`include "carryLookahead16.v"
module fastAdder2Stage(
    input clock,
    input reset,
    input [31:0] in_a,
    input [31:0] in_b,
    output [32:0] out_sum
);

parameter WIDTH = 32;

// buffer registers for IO
reg [WIDTH-1:0] buffer_in_a;
reg [WIDTH-1:0] buffer_in_b;
reg [WIDTH:0] buffer_out_sum;

// stage 1 pipeline registers
reg [(WIDTH/2 -1):0] pipeline_in_a;   //for higher 16 bits of in_a
reg [(WIDTH/2 -1):0] pipeline_in_b;   //for higher 16 bits of in_b
reg [(WIDTH/2):0] pipeline_sum0;   //for {carry,sum} generated by adder0


// wire fot stage 1 output --- carry is the MSB bit
wire [(WIDTH/2):0] sum0;

CLA_16bit cla0(
    buffer_in_a[(WIDTH/2 - 1):0],
    buffer_in_b[(WIDTH/2 - 1):0],
    1'b0,
    sum0[(WIDTH/2 - 1):0],
    sum0[(WIDTH/2)]);

always @(posedge clock) begin
    if (reset) begin
        pipeline_in_a <= {(WIDTH/2 - 1){1'b0}};
        pipeline_in_b <= {(WIDTH/2 - 1){1'b0}};
        pipeline_sum0 <= {(WIDTH/2){1'b0}};
    end 
    else begin
        buffer_in_a <= in_a;
        buffer_in_b <= in_b;

        pipeline_in_a <= buffer_in_a[(WIDTH-1):(WIDTH/2)];
        pipeline_in_b <= buffer_in_b[(WIDTH-1):(WIDTH/2)];

        pipeline_sum0 <= sum0;        
    end    
end

// stage 2
wire [(WIDTH/2):0] sum1;

CLA_16bit cla1(
    pipeline_in_a,
    pipeline_in_b,
    sum0[(WIDTH/2)],
    sum1[(WIDTH/2 - 1):0],
    sum1[(WIDTH/2)]
);

always @(posedge clock) begin
    if (reset) begin
        // flush output buffer
        buffer_out_sum <= {WIDTH{1'b0}};
    end 
    else begin
        buffer_out_sum <= {sum1, pipeline_sum0};
    end
end

assign out_sum = buffer_out_sum;
    
endmodule