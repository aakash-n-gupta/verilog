// result shows 0 if bits are unequal an 1 only when both x and y are equal

module comparator (
    parameter WIDTH = 8;

    input x[WIDTH - 1:0],
    input y{WIDTH - 1:0},
    output result
);

    assign 
    
endmodule