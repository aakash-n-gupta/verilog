module adderGenerator #(parameter WIDTH = 16) (
    input [WIDTH -1 : 0] in_a, 
    input [WIDTH -1 : 0] in_b, 
    input in_carry,
    output [WIDTH - 1 : 0] sum,
    output out_carry 
    );
    assign {out_carry, sum} = in_a + in_b + in_carry;
endmodule

module adder2StageBuf (
    input clock,
    input reset,
    input[31:0] in_a,
    input[31:0] in_b,
    output[32:0] out_sum    // 32 bit sum is easier to debug in simulation
    // output out_carry -- //use for synthesys, 
);

    parameter WIDTH = 32;
    
    // buffer registers for IO ports
    reg [WIDTH-1:0] buffer_in_a;
    reg [WIDTH-1:0] buffer_in_b;
    reg [WIDTH:0] buffer_out_sum;

    // stage 1 pipeline registers
    reg [(WIDTH/2 -1):0] pipeline_in_a;   //for higher 16 bits of in_a
    reg [(WIDTH/2 -1):0] pipeline_in_b;   //for higher 16 bits of in_b
    reg [(WIDTH/2 -1):0] pipeline_sum0;   //for sum generated by adder0
    reg pipeline_carry0;        //for carry_out generated by adder0

    // wires for stage 1 outputs
    wire [(WIDTH/2 -1):0] sum0;
    wire carry0;

    // carryin for adder0 is set to 0.
    // sending the output directly to the pipeline regs, no explicit wires declared
    adderGenerator adder0(buffer_in_a[15:0], buffer_in_b[15:0], 1'b0, sum0, carry0);

    always @(posedge clock) begin
        if(reset)
        begin
            // resets all pipeline_regs of stage 1 to 0
            pipeline_in_a <= {(WIDTH/2 - 1){1'b0}};
            pipeline_in_b <= {(WIDTH/2 - 1){1'b0}};
            pipeline_sum0 <= {(WIDTH/2 - 1){1'b0}};
            pipeline_carry0 <= 1'b0;
        end
        else begin
            // buffer IO stage
            buffer_in_a <= in_a;
            buffer_in_b <= in_b;

            pipeline_in_a <= buffer_in_a[(WIDTH-1):(WIDTH/2)];
            pipeline_in_b <= buffer_in_b[(WIDTH-1):(WIDTH/2)];

            pipeline_sum0 <= sum0;
            pipeline_carry0 <= carry0;            
        end
        
    end

    // wires for stage 2 output
    wire [(WIDTH/2 - 1):0] sum1;
    wire carry1;

    adderGenerator adder1 (pipeline_in_a, pipeline_in_b, pipeline_carry0, sum1[(WIDTH/2 - 1):0], carry1);

    always @(posedge clock ) begin
        if (reset) begin
            // flush output buffer
            buffer_out_sum <= {(WIDTH+1){1'b0}};
        end
        else begin
            buffer_out_sum <= {carry1, sum1 ,pipeline_sum0};
        end
        
    end

    assign out_sum = buffer_out_sum;


endmodule