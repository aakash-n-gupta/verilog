module carryLookaheadFA (
    input in_a,
    input in_b,
    input in_carry,
    output out_sum,
    output out_carry
);
    wire propogate;
    wire lookahead;

    assign out_sum = 
endmodule